
module c10_clkctrl (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
